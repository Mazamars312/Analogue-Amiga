module amiga_keyboard_convert (
input clk,
input [7:0] input_keyboard,
output reg [7:0] output_keyboard
);

reg [7:0] mem [255:0];

initial begin
mem[0  ] <=	8'h00;            /**< 0   KEY_RESERVED */
mem[1  ] <=	8'h45;              /**< 1   KEY_ESC */
mem[2  ] <=	8'h01;              /**< 2   KEY_1 */
mem[3  ] <=	8'h02;              /**< 3   KEY_2 */
mem[4  ] <=	8'h03;              /**< 4   KEY_3 */
mem[5  ] <=	8'h04;              /**< 5   KEY_4 */
mem[6  ] <=	8'h05;              /**< 6   KEY_5 */
mem[7  ] <=	8'h06;              /**< 7   KEY_6 */
mem[8  ] <=	8'h07;              /**< 8   KEY_7 */
mem[9  ] <=	8'h08;              /**< 9   KEY_8 */
mem[10 ] <=	8'h09;              /**< 10  KEY_9 */
mem[11 ] <=	8'h0a;              /**< 11  KEY_0 */
mem[12 ] <=	8'h0b;              /**< 12  KEY_MINUS */
mem[13 ] <=	8'h0c;              /**< 13  KEY_EQUAL */
mem[14 ] <=	8'h41;              /**< 14  KEY_BACKSPACE */
mem[15 ] <=	8'h42;              /**< 15  KEY_TAB */
mem[16 ] <=	8'h10;              /**< 16  KEY_Q */
mem[17 ] <=	8'h11;              /**< 17  KEY_W */
mem[18 ] <=	8'h12;              /**< 18  KEY_E */
mem[19 ] <=	8'h13;              /**< 19  KEY_R */
mem[20 ] <=	8'h14;              /**< 20  KEY_T */
mem[21 ] <=	8'h15;              /**< 21  KEY_Y */
mem[22 ] <=	8'h16;              /**< 22  KEY_U */
mem[23 ] <=	8'h17;              /**< 23  KEY_I */
mem[24 ] <=	8'h18;              /**< 24  KEY_O */
mem[25 ] <=	8'h19;              /**< 25  KEY_P */
mem[26 ] <=	8'h1a;              /**< 26  KEY_LEFTBRACE */
mem[27 ] <=	8'h1b;              /**< 27  KEY_RIGHTBRACE */
mem[28 ] <=	8'h44;              /**< 28  KEY_ENTER */
mem[29 ] <=	8'h63;              /**< 29  KEY_LEFTCTRL */
mem[30 ] <=	8'h20;              /**< 30  KEY_A */
mem[31 ] <=	8'h21;              /**< 31  KEY_S */
mem[32 ] <=	8'h22;              /**< 32  KEY_D */
mem[33 ] <=	8'h23;              /**< 33  KEY_F */
mem[34 ] <=	8'h24;              /**< 34  KEY_G */
mem[35 ] <=	8'h25;              /**< 35  KEY_H */
mem[36 ] <=	8'h26;              /**< 36  KEY_J */
mem[37 ] <=	8'h27;              /**< 37  KEY_K */
mem[38 ] <=	8'h28;              /**< 38  KEY_L */
mem[39 ] <=	8'h29;              /**< 39  KEY_SEMICOLON */
mem[40 ] <=	8'h2a;              /**< 40  KEY_APOSTROPHE */
mem[41 ] <=	8'h00;              /**< 41  KEY_GRAVE */
mem[42 ] <=	8'h60;              /**< 42  KEY_LEFTSHIFT */
mem[43 ] <=	8'h0d;              /**< 43  KEY_BACKSLASH */
mem[44 ] <=	8'h31;              /**< 44  KEY_Z */
mem[45 ] <=	8'h32;              /**< 45  KEY_X */
mem[46 ] <=	8'h33;              /**< 46  KEY_C */
mem[47 ] <=	8'h34;              /**< 47  KEY_V */
mem[48 ] <=	8'h35;              /**< 48  KEY_B */
mem[49 ] <=	8'h36;              /**< 49  KEY_N */
mem[50 ] <=	8'h37;              /**< 50  KEY_M */
mem[51 ] <=	8'h38;              /**< 51  KEY_COMMA */
mem[52 ] <=	8'h39;              /**< 52  KEY_DOT */
mem[53 ] <=	8'h3a;              /**< 53  KEY_SLASH */
mem[54 ] <=	8'h61;              /**< 54  KEY_RIGHTSHIFT */
mem[55 ] <=	8'h5d;              /**< 55  KEY_KPASTERISK */
mem[56 ] <=	8'h64;              /**< 56  KEY_LEFTALT */
mem[57 ] <=	8'h40;              /**< 57  KEY_SPACE */
mem[58 ] <=	8'h62;/**< 58  KEY_CAPSLOCK */
mem[59 ] <=	8'h50;              /**< 59  KEY_F1 */
mem[60 ] <=	8'h51;              /**< 60  KEY_F2 */
mem[61 ] <=	8'h52;              /**< 61  KEY_F3 */
mem[62 ] <=	8'h53;              /**< 62  KEY_F4 */
mem[63 ] <=	8'h54;              /**< 63  KEY_F5 */
mem[64 ] <=	8'h55;              /**< 64  KEY_F6 */
mem[65 ] <=	8'h56;              /**< 65  KEY_F7 */
mem[66 ] <=	8'h57;              /**< 66  KEY_F8 */
mem[67 ] <=	8'h58;              /**< 67  KEY_F9 */
mem[68 ] <=	8'h59;              /**< 68  KEY_F10 */
mem[69 ] <=	8'h00;            /**< 69  KEY_NUMLOCK */
mem[70 ] <=	8'h00;            /**< 70  KEY_SCROLLLOCK */
mem[71 ] <=	8'h3d;              /**< 71  KEY_KP7 */
mem[72 ] <=	8'h3e;              /**< 72  KEY_KP8 */
mem[73 ] <=	8'h3f;              /**< 73  KEY_KP9 */
mem[74 ] <=	8'h4a;              /**< 74  KEY_KPMINUS */
mem[75 ] <=	8'h2d;              /**< 75  KEY_KP4 */
mem[76 ] <=	8'h2e;              /**< 76  KEY_KP5 */
mem[77 ] <=	8'h2f;              /**< 77  KEY_KP6 */
mem[78 ] <=	8'h5e;              /**< 78  KEY_KPPLUS */
mem[79 ] <=	8'h1d;              /**< 79  KEY_KP1 */
mem[80 ] <=	8'h1e;              /**< 80  KEY_KP2 */
mem[81 ] <=	8'h1f;              /**< 81  KEY_KP3 */
mem[82 ] <=	8'h0f;              /**< 82  KEY_KP0 */
mem[83 ] <=	8'h3c;              /**< 83  KEY_KPDOT */
mem[84 ] <=	8'h00;            /**< 84  ??? */
mem[85 ] <=	8'h00;            /**< 85  KEY_ZENKAKU */
mem[86 ] <=	8'h30;              /**< 86  KEY_102ND; '<' on most keyboards */
mem[87 ] <=	8'h5f;              /**< 87  KEY_F11 */
mem[88 ] <=	8'h00;            /**< 88  KEY_F12 */
mem[89 ] <=	8'h00;            /**< 89  KEY_RO */
mem[90 ] <=	8'h00;            /**< 90  KEY_KATAKANA */
mem[91 ] <=	8'h00;            /**< 91  KEY_HIRAGANA */
mem[92 ] <=	8'h00;            /**< 92  KEY_HENKAN */
mem[93 ] <=	8'h00;            /**< 93  KEY_KATAKANA */
mem[94 ] <=	8'h00;            /**< 94  KEY_MUHENKAN */
mem[95 ] <=	8'h00;            /**< 95  KEY_KPJPCOMMA */
mem[96 ] <=	8'h43;              /**< 96  KEY_KPENTER */
mem[97 ] <=	8'h63;              /**< 97  KEY_RIGHTCTRL */
mem[98 ] <=	8'h5c;              /**< 98  KEY_KPSLASH */
mem[99 ] <=	8'h00;            /**< 99  KEY_SYSRQ */
mem[100] <=	8'h65;              /**< 100 KEY_RIGHTALT */
mem[101] <=	8'h00;            /**< 101 KEY_LINEFEED */
mem[102] <=	8'h6a;              /**< 102 KEY_HOME */
mem[103] <=	8'h4c;              /**< 103 KEY_UP */
mem[104] <=	8'h5b;              /**< 104 KEY_PAGEUP */
mem[105] <=	8'h4f;              /**< 105 KEY_LEFT */
mem[106] <=	8'h4e;              /**< 106 KEY_RIGHT */
mem[107] <=	8'h00;            /**< 107 KEY_END */
mem[108] <=	8'h4d;              /**< 108 KEY_DOWN */
mem[109] <=	8'h5a;              /**< 109 KEY_PAGEDOWN */
mem[110] <=	8'h0d;              /**< 110 KEY_INSERT */
mem[111] <=	8'h46;              /**< 111 KEY_DELETE */
mem[112] <=	8'h00;            /**< 112 KEY_MACRO */
mem[113] <=	8'h00;            /**< 113 KEY_MUTE */
mem[114] <=	8'h00;            /**< 114 KEY_VOLUMEDOWN */
mem[115] <=	8'h00;            /**< 115 KEY_VOLUMEUP */
mem[116] <=	8'h00;            /**< 116 KEY_POWER */
mem[117] <=	8'h00;            /**< 117 KEY_KPEQUAL */
mem[118] <=	8'h00;            /**< 118 KEY_KPPLUSMINUS */
mem[119] <=	8'h00;            /**< 119 KEY_PAUSE */
mem[120] <=	8'h00;            /**< 120 KEY_SCALE */
mem[121] <=	8'h00;            /**< 121 KEY_KPCOMMA */
mem[122] <=	8'h00;            /**< 122 KEY_HANGEUL */
mem[123] <=	8'h00;            /**< 123 KEY_HANJA */
mem[124] <=	8'h00;            /**< 124 KEY_YEN */
mem[125] <=	8'h66;              /**< 125 KEY_LEFTMETA */
mem[126] <=	8'h67;              /**< 126 KEY_RIGHTMETA */
mem[127] <=	8'h00;            /**< 127 KEY_COMPOSE */
mem[128] <=	8'h00;            /**< 128 KEY_STOP */
mem[129] <=	8'h00;            /**< 129 KEY_AGAIN */
mem[130] <=	8'h00;            /**< 130 KEY_PROPS */
mem[131] <=	8'h00;            /**< 131 KEY_UNDO */
mem[132] <=	8'h00;            /**< 132 KEY_FRONT */
mem[133] <=	8'h00;            /**< 133 KEY_COPY */
mem[134] <=	8'h00;            /**< 134 KEY_OPEN */
mem[135] <=	8'h00;            /**< 135 KEY_PASTE */
mem[136] <=	8'h00;            /**< 136 KEY_FIND */
mem[137] <=	8'h00;            /**< 137 KEY_CUT */
mem[138] <=	8'h00;            /**< 138 KEY_HELP */
mem[139] <=	8'h00;            /**< 139 KEY_MENU */
mem[140] <=	8'h00;            /**< 140 KEY_CALC */
mem[141] <=	8'h00;            /**< 141 KEY_SETUP */
mem[142] <=	8'h00;            /**< 142 KEY_SLEEP */
mem[143] <=	8'h00;            /**< 143 KEY_WAKEUP */
mem[144] <=	8'h00;            /**< 144 KEY_FILE */
mem[145] <=	8'h00;            /**< 145 KEY_SENDFILE */
mem[146] <=	8'h00;            /**< 146 KEY_DELETEFILE */
mem[147] <=	8'h00;            /**< 147 KEY_XFER */
mem[148] <=	8'h00;            /**< 148 KEY_PROG1 */
mem[149] <=	8'h00;            /**< 149 KEY_PROG2 */
mem[150] <=	8'h00;            /**< 150 KEY_WWW */
mem[151] <=	8'h00;            /**< 151 KEY_MSDOS */
mem[152] <=	8'h00;            /**< 152 KEY_SCREENLOCK */
mem[153] <=	8'h00;            /**< 153 KEY_DIRECTION */
mem[154] <=	8'h00;            /**< 154 KEY_CYCLEWINDOWS */
mem[155] <=	8'h00;            /**< 155 KEY_MAIL */
mem[156] <=	8'h00;            /**< 156 KEY_BOOKMARKS */
mem[157] <=	8'h00;            /**< 157 KEY_COMPUTER */
mem[158] <=	8'h00;            /**< 158 KEY_BACK */
mem[159] <=	8'h00;            /**< 159 KEY_FORWARD */
mem[160] <=	8'h00;            /**< 160 KEY_CLOSECD */
mem[161] <=	8'h00;            /**< 161 KEY_EJECTCD */
mem[162] <=	8'h00;            /**< 162 KEY_EJECTCLOSECD */
mem[163] <=	8'h00;            /**< 163 KEY_NEXTSONG */
mem[164] <=	8'h00;            /**< 164 KEY_PLAYPAUSE */
mem[165] <=	8'h00;            /**< 165 KEY_PREVIOUSSONG */
mem[166] <=	8'h00;            /**< 166 KEY_STOPCD */
mem[167] <=	8'h00;            /**< 167 KEY_RECORD */
mem[168] <=	8'h00;            /**< 168 KEY_REWIND */
mem[169] <=	8'h00;            /**< 169 KEY_PHONE */
mem[170] <=	8'h00;            /**< 170 KEY_ISO */
mem[171] <=	8'h00;            /**< 171 KEY_CONFIG */
mem[172] <=	8'h00;            /**< 172 KEY_HOMEPAGE */
mem[173] <=	8'h00;            /**< 173 KEY_REFRESH */
mem[174] <=	8'h00;            /**< 174 KEY_EXIT */
mem[175] <=	8'h00;            /**< 175 KEY_MOVE */
mem[176] <=	8'h00;            /**< 176 KEY_EDIT */
mem[177] <=	8'h00;            /**< 177 KEY_SCROLLUP */
mem[178] <=	8'h00;            /**< 178 KEY_SCROLLDOWN */
mem[179] <=	8'h00;            /**< 179 KEY_KPLEFTPAREN */
mem[180] <=	8'h00;            /**< 180 KEY_KPRIGHTPAREN */
mem[181] <=	8'h00;            /**< 181 KEY_NEW */
mem[182] <=	8'h00;            /**< 182 KEY_REDO */
mem[183] <=	8'h5a;              /**< 183 KEY_F13 */
mem[184] <=	8'h5b;              /**< 184 KEY_F14 */
mem[185] <=	8'h00;            /**< 185 KEY_F15 */
mem[186] <=	8'h5f;              /**< 186 KEY_F16 */
mem[187] <=	8'h00;            /**< 187 KEY_F17 */
mem[188] <=	8'h00;            /**< 188 KEY_F18 */
mem[189] <=	8'h00;            /**< 189 KEY_F19 */
mem[190] <=	8'h00;            /**< 190 KEY_F20 */
mem[191] <=	8'h00;            /**< 191 KEY_F21 */
mem[192] <=	8'h00;            /**< 192 KEY_F22 */
mem[193] <=	8'h00;            /**< 193 KEY_F23 */
mem[194] <=	8'h2b;              /**< 194 # on German keyboard; was 8'h63 (CTRL on Amiga); 194 KEY_F24 */
mem[195] <=	8'h00;            /**< 195 ??? */
mem[196] <=	8'h00;            /**< 196 ??? */
mem[197] <=	8'h00;            /**< 197 ??? */
mem[198] <=	8'h00;            /**< 198 ??? */
mem[199] <=	8'h00;            /**< 199 ??? */
mem[200] <=	8'h00;            /**< 200 KEY_PLAYCD */
mem[201] <=	8'h00;            /**< 201 KEY_PAUSECD */
mem[202] <=	8'h00;            /**< 202 KEY_PROG3 */
mem[203] <=	8'h00;            /**< 203 KEY_PROG4 */
mem[204] <=	8'h00;            /**< 204 KEY_DASHBOARD */
mem[205] <=	8'h00;            /**< 205 KEY_SUSPEND */
mem[206] <=	8'h00;            /**< 206 KEY_CLOSE */
mem[207] <=	8'h00;            /**< 207 KEY_PLAY */
mem[208] <=	8'h00;            /**< 208 KEY_FASTFORWARD */
mem[209] <=	8'h00;            /**< 209 KEY_BASSBOOST */
mem[210] <=	8'h00;            /**< 210 KEY_PRINT */
mem[211] <=	8'h00;            /**< 211 KEY_HP */
mem[212] <=	8'h00;            /**< 212 KEY_CAMERA */
mem[213] <=	8'h00;            /**< 213 KEY_SOUND */
mem[214] <=	8'h00;            /**< 214 KEY_QUESTION */
mem[215] <=	8'h00;            /**< 215 KEY_EMAIL */
mem[216] <=	8'h00;            /**< 216 KEY_CHAT */
mem[217] <=	8'h00;            /**< 217 KEY_SEARCH */
mem[218] <=	8'h00;            /**< 218 KEY_CONNECT */
mem[219] <=	8'h00;            /**< 219 KEY_FINANCE */
mem[220] <=	8'h00;            /**< 220 KEY_SPORT */
mem[221] <=	8'h00;            /**< 221 KEY_SHOP */
mem[222] <=	8'h00;            /**< 222 KEY_ALTERASE */
mem[223] <=	8'h00;            /**< 223 KEY_CANCEL */
mem[224] <=	8'h00;            /**< 224 KEY_BRIGHT_DOWN */
mem[225] <=	8'h00;            /**< 225 KEY_BRIGHT_UP */
mem[226] <=	8'h00;            /**< 226 KEY_MEDIA */
mem[227] <=	8'h00;            /**< 227 KEY_SWITCHVIDEO */
mem[228] <=	8'h00;            /**< 228 KEY_DILLUMTOGGLE */
mem[229] <=	8'h00;            /**< 229 KEY_DILLUMDOWN */
mem[230] <=	8'h00;            /**< 230 KEY_DILLUMUP */
mem[231] <=	8'h00;            /**< 231 KEY_SEND */
mem[232] <=	8'h00;            /**< 232 KEY_REPLY */
mem[233] <=	8'h00;            /**< 233 KEY_FORWARDMAIL */
mem[234] <=	8'h00;            /**< 234 KEY_SAVE */
mem[235] <=	8'h00;            /**< 235 KEY_DOCUMENTS */
mem[236] <=	8'h00;            /**< 236 KEY_BATTERY */
mem[237] <=	8'h00;            /**< 237 KEY_BLUETOOTH */
mem[238] <=	8'h00;            /**< 238 KEY_WLAN */
mem[239] <=	8'h00;            /**< 239 KEY_UWB */
mem[240] <=	8'h00;            /**< 240 KEY_UNKNOWN */
mem[241] <=	8'h00;            /**< 241 KEY_VIDEO_NEXT */
mem[242] <=	8'h00;            /**< 242 KEY_VIDEO_PREV */
mem[243] <=	8'h00;            /**< 243 KEY_BRIGHT_CYCLE */
mem[244] <=	8'h00;            /**< 244 KEY_BRIGHT_AUTO */
mem[245] <=	8'h00;            /**< 245 KEY_DISPLAY_OFF */
mem[246] <=	8'h00;            /**< 246 KEY_WWAN */
mem[247] <=	8'h00;            /**< 247 KEY_RFKILL */
mem[248] <=	8'h00;            /**< 248 KEY_MICMUTE */
mem[249] <=	8'h00;            /**< 249 ??? */
mem[250] <=	8'h00;            /**< 250 ??? */
mem[251] <=	8'h00;            /**< 251 ??? */
mem[252] <=	8'h00;            /**< 252 ??? */
mem[253] <=	8'h00;            /**< 253 ??? */
mem[254] <=	8'h00;            /**< 254 ??? */
mem[255] <=	8'h00;            /**< 255 ??? */

end


always @(posedge clk) output_keyboard <= mem[input_keyboard];


endmodule